library verilog;
use verilog.vl_types.all;
entity main_AES_vlg_vec_tst is
end main_AES_vlg_vec_tst;
