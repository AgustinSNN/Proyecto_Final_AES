library verilog;
use verilog.vl_types.all;
entity key_expansion_vlg_vec_tst is
end key_expansion_vlg_vec_tst;
